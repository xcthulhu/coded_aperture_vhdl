../vhdl/common_decs.vhdl