../vhdl/rstgen_syscon.vhdl