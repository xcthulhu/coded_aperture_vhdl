../vhdl/top_mod.vhdl