../vhdl/wb_fifo_chain.vhdl