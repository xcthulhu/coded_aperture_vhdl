../vhdl/sclk_data_acq.vhdl