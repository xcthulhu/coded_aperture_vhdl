Library c;
Use c.stdio_h.all;

Entity hello is
End Entity hello;

Architecture test of hello is
Begin
  printf("Hello World!\n");
End Architecture test;
