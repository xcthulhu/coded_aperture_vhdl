../vhdl/intercon.vhdl