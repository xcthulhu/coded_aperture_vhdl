../vhdl/wishbone_wrapper.vhdl