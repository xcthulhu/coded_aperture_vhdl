../vhdl/irq_mngr.vhdl