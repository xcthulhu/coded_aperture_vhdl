../vhdl/intercon_decs.vhdl