../vhdl/wb_fifo.vhdl