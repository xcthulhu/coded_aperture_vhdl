../vhdl/data_bridge.vhdl