../vhdl/fifo.vhdl